//-------------------------------------------------------------------------
//      VGA controller                                                   --
//      Kyle Kloepper                                                    --
//      4-05-2005                                                        --
//                                                                       --
//      Modified by Stephen Kempf 04-08-2005                             --
//                                10-05-2006                             --
//                                03-12-2007                             --
//      Translated by Joe Meng    07-07-2013                             --
//      Modified by Po-Han Huang  12-08-2017                             --
//      Spring 2018 Distribution                                         --
//                                                                       --
//      Used standard 640x480 vga found at epanorama                     --
//                                                                       --
//      reference: http://www.xilinx.com/bvdocs/userguides/ug130.pdf     --
//                 http://www.epanorama.net/documents/pc/vga_timing.html --
//                                                                       --
//      note: The standard is changed slightly because of 25 mhz instead --
//            of 25.175 mhz pixel clock. Refresh rate drops slightly.    --
//                                                                       --
//      For use with ECE 385 Lab 8 and Final Project                     --
//      ECE Department @ UIUC                                            --
//-------------------------------------------------------------------------


module  VGA_controller (input              Clk,         // 50 MHz clock
                                           Reset,       // Active-high reset signal
                        output logic       VGA_HS,      // Horizontal sync pulse.  Active low
                                           VGA_VS,      // Vertical sync pulse.  Active low
                        input              VGA_CLK,     // 25 MHz VGA clock input
                        output logic       VGA_BLANK_N, // Blanking interval indicator.  Active low.
                                           VGA_SYNC_N,  // Composite Sync signal.  Active low.  We don't use it in this lab,
                                                        // but the video DAC on the DE2 board requires an input for it.
                        output logic [9:0] DrawX,       // horizontal coordinate
                                           DrawY        // vertical coordinate
                        );     
    
    // 800 pixels per line (including front/back porch)
    // 525 lines per frame (including front/back porch)
    parameter [9:0] H_TOTAL = 10'd800;
    parameter [9:0] V_TOTAL = 10'd525;
    
    logic VGA_HS_in, VGA_VS_in, VGA_BLANK_N_in;
    logic [9:0] h_counter, v_counter;
    logic [9:0] h_counter_in, v_counter_in;
    
    assign VGA_SYNC_N = 1'b0;
    assign DrawX = h_counter;
    assign DrawY = v_counter;
    
    // VGA control signals. 
    // VGA_CLK is generated by PLL, so you will have to manually generate it in simulation.
    always_ff @ (posedge VGA_CLK)
    begin
        if (Reset)
        begin
            VGA_HS <= 1'b0;
            VGA_VS <= 1'b0;
            VGA_BLANK_N <= 1'b0;
            h_counter <= 10'd0;
            v_counter <= 10'd0;
        end
        else
        begin
            VGA_HS <= VGA_HS_in;
            VGA_VS <= VGA_VS_in;
            VGA_BLANK_N <= VGA_BLANK_N_in;
            h_counter <= h_counter_in;
            v_counter <= v_counter_in;
        end
    end
    
    always_comb
    begin
        // horizontal and vertical counter
        h_counter_in = h_counter + 10'd1;
        v_counter_in = v_counter;
        if(h_counter + 10'd1 == H_TOTAL)
        begin
            h_counter_in = 10'd0;
            if(v_counter + 10'd1 == V_TOTAL)
                v_counter_in = 10'd0;
            else
                v_counter_in = v_counter + 10'd1;
        end
        // Horizontal sync pulse is 96 pixels long at pixels 656-752
        // (Signal is registered to ensure clean output waveform)
        VGA_HS_in = 1'b1;
        if(h_counter_in >= 10'd656 && h_counter_in < 10'd752)
            VGA_HS_in = 1'b0;
        // Vertical sync pulse is 2 lines (800 pixels each) long at line 490-491
        //(Signal is registered to ensure clean output waveform)
        VGA_VS_in = 1'b1;
        if(v_counter_in >= 10'd490 && v_counter_in < 10'd492)
            VGA_VS_in = 1'b0;
        // Display pixels (inhibit blanking) between horizontal 0-639 and vertical 0-479 (640x480)
        VGA_BLANK_N_in = 1'b0;
        if(h_counter_in < 10'd640 && v_counter_in < 10'd480)
            VGA_BLANK_N_in = 1'b1;
    end
    
endmodule


module VGA_mapper(
    input logic CLK, VGA_CLK, RESET,
    input logic [1:0] VGA_ADDR,
    input logic [31:0] VGA_WRITEDATA,
    output logic [31:0] VGA_READDATA,
    input logic [3:0] VGA_BYTE_EN,
    input logic VGA_WRITE, VGA_CS, VGA_READ,
    input logic VGA_BLANK_N,
    output logic [7:0] VGA_R, VGA_G, VGA_B,

    // Avalon-MM Master Signals
    output logic [31:0] VGA_MASTER_ADDR,
    output logic VGA_MASTER_READ,
    input  logic [31:0] VGA_MASTER_READDATA,
    output logic VGA_MASTER_CS,
    input  logic VGA_MASTER_WAIT_REQUEST,
    input logic  VGA_MASTER_READDATAVALID,

    input logic [9:0] DrawX,
    input logic [9:0] DrawY,

    output logic [7:0] DEBUG

);

    logic [31:0] ram1_data, ram2_data;
    logic ram1_we, ram2_we;
    logic current_ram = 0;

    logic [31:0] copy_counter = 0, copy_counter_next; // coping offset from start of line
    logic [31:0] offset_counter = 0, offset_counter_next; // num lines offset from start

    logic [31:0] frame_pointer = 0, frame_pointer_next; // location of image 
    logic [31:0] should_draw = 0, should_draw_next; // TODO

     enum logic [3:0] {
             IDLE,
             COPYING,
             COPYING1,
             COPYING2,
             COPYING3,
             COPYING4
         }   State, Next_state; // Data Copy State

    
    vga_ram #(0) ram1(.output_data(ram1_data),
        .input_data(VGA_MASTER_READDATA), 
        .write_address(copy_counter), .read_address(DrawX),
        .we(ram1_we), .clk(CLK), .read_clk(VGA_CLK));

    vga_ram #(1) ram2(.output_data(ram2_data),
        .input_data(VGA_MASTER_READDATA), 
        .write_address(copy_counter), .read_address(DrawX),
        .we(ram2_we), .clk(CLK), .read_clk(VGA_CLK));


    always_comb begin
        DEBUG = 1;
        frame_pointer_next = frame_pointer;
        should_draw_next = should_draw;
        copy_counter_next = copy_counter;
        offset_counter_next = offset_counter;
        VGA_READDATA = 4'hzzzz;
        ram1_we = 0;
        ram2_we = 0;

        // Master default values
        VGA_MASTER_ADDR = 4'hzzzz;
        VGA_MASTER_CS = 0;
        VGA_MASTER_READ = 0;

        // Slave read writes
        if(VGA_CS) begin
            if(VGA_WRITE) begin
                if(VGA_ADDR == 0) 
                    frame_pointer_next = VGA_WRITEDATA;
                if(VGA_ADDR == 1) 
                    should_draw_next = VGA_WRITEDATA;
            end else if(VGA_READ) begin
                if(VGA_ADDR == 0) 
                    VGA_READDATA = frame_pointer;
                if(VGA_ADDR == 1) 
                    VGA_READDATA = should_draw;
            end
        end

        if(~(State == IDLE)) begin
           // ram1_we = (current_ram == 1); // Write to R1 if reading from R2
           // ram2_we = (current_ram == 0); // Write to R2 if reading from R1
            ram1_we = 1;
            VGA_MASTER_CS = 1;
            VGA_MASTER_READ = 1;
            VGA_MASTER_ADDR = frame_pointer + ((640*(DrawY))+copy_counter) * 4;
        end
        //VGA_MASTER_ADDR = frame_pointer + ((640*DrawY)+DrawX) * 4;

        unique case (State)
            IDLE: begin
                if((DrawX <= 640) & (DrawY <= 480))
                    Next_state = COPYING;
                else begin
                    Next_state = IDLE;
                    if (DrawY > 480)
                        offset_counter_next = 0;
                end
            end
            COPYING: begin
                //if(VGA_MASTER_WAIT_REQUEST)
                //    Next_state = COPYING;
                //else 
                if (copy_counter == 639) begin
                    Next_state = IDLE;
                    copy_counter_next = 0;
                    offset_counter_next = offset_counter + 1;
                end else begin
                    //if (VGA_MASTER_READDATAVALID) begin
                    if (~VGA_MASTER_WAIT_REQUEST) begin
                        Next_state = COPYING1;
                    end else begin
                        Next_state = COPYING;
                    end
                end
            end
            COPYING1: begin
                    Next_state = COPYING;
                    copy_counter_next = copy_counter + 1;
            end
            default:
                Next_state = State;
        endcase
    end

    // D flop flops
    always_ff @(posedge CLK) begin //50 MHz
        if (RESET) begin
            frame_pointer <= 0;
            should_draw <= 0;
            State <= IDLE;
            copy_counter <= 0;
            offset_counter <= 0;
        end else begin
            frame_pointer <= frame_pointer_next;
            should_draw <= should_draw_next;
            State <= Next_state;
            copy_counter <= copy_counter_next;
            offset_counter <= offset_counter_next;
        end
    end

     always_ff @(posedge VGA_CLK) begin // 25 MHz

             //VGA_R <= VGA_MASTER_READDATA[7:0];
             //VGA_G <= VGA_MASTER_READDATA[15:8];
             //VGA_B <= VGA_MASTER_READDATA[23:16];
             VGA_R <= ram1_data[7:0];
             VGA_G <= ram1_data[15:8];
             VGA_B <= ram1_data[23:16];
 
//         if(current_ram == 0) begin
//             VGA_R <= ram1_data[7:0];
//             VGA_G <= ram1_data[15:8];
//             VGA_B <= ram1_data[23:16];
//         end else begin
//             VGA_R <= ram1_data[7:0];
//             VGA_G <= ram1_data[15:8];
//             VGA_B <= ram1_data[23:16];
//         end
 
 
     end
     
 
endmodule

module vga_ram #(parameter ram_num = 0)(
    output logic [31:0] output_data,
    input logic [31:0] input_data,
    input [10:0] write_address, read_address,
    input we, clk, read_clk
);

logic [31:0] mem[640];

initial
begin
    if(ram_num == 0) begin
        $display("Reading ram 0");
        $readmemh("vga_ram0.txt", mem);
    end else if(ram_num == 1) begin
        $display("Reading ram 1");
        $readmemh("vga_ram1.txt", mem);
    end else begin
        $display("Unknown ram number----------------------");
    end
end

always_ff @ (posedge clk) begin
    if (we)
        mem[write_address] <= input_data;
end

always_ff @ (posedge read_clk) begin
    output_data <= mem[read_address];
end
endmodule
