//-------------------------------------------------------------------------
//      VGA controller                                                   --
//      Kyle Kloepper                                                    --
//      4-05-2005                                                        --
//                                                                       --
//      Modified by Stephen Kempf 04-08-2005                             --
//                                10-05-2006                             --
//                                03-12-2007                             --
//      Translated by Joe Meng    07-07-2013                             --
//      Modified by Po-Han Huang  12-08-2017                             --
//      Spring 2018 Distribution                                         --
//                                                                       --
//      Used standard 640x480 vga found at epanorama                     --
//                                                                       --
//      reference: http://www.xilinx.com/bvdocs/userguides/ug130.pdf     --
//                 http://www.epanorama.net/documents/pc/vga_timing.html --
//                                                                       --
//      note: The standard is changed slightly because of 25 mhz instead --
//            of 25.175 mhz pixel clock. Refresh rate drops slightly.    --
//                                                                       --
//      For use with ECE 385 Lab 8 and Final Project                     --
//      ECE Department @ UIUC                                            --
//-------------------------------------------------------------------------


module  VGA_controller (input              Clk,         // 50 MHz clock
                                           Reset,       // Active-high reset signal
                        output logic       VGA_HS,      // Horizontal sync pulse.  Active low
                                           VGA_VS,      // Vertical sync pulse.  Active low
                        input              VGA_CLK,     // 25 MHz VGA clock input
                        output logic       VGA_BLANK_N, // Blanking interval indicator.  Active low.
                                           VGA_SYNC_N,  // Composite Sync signal.  Active low.  We don't use it in this lab,
                                                        // but the video DAC on the DE2 board requires an input for it.
                        output logic [9:0] DrawX,       // horizontal coordinate
                                           DrawY        // vertical coordinate
                        );     
    
    // 800 pixels per line (including front/back porch)
    // 525 lines per frame (including front/back porch)
    parameter [9:0] H_TOTAL = 10'd800;
    parameter [9:0] V_TOTAL = 10'd525;
    
    logic VGA_HS_in, VGA_VS_in, VGA_BLANK_N_in;
    logic [9:0] h_counter, v_counter;
    logic [9:0] h_counter_in, v_counter_in;
    
    assign VGA_SYNC_N = 1'b0;
    assign DrawX = h_counter;
    assign DrawY = v_counter;
    
    // VGA control signals. 
    // VGA_CLK is generated by PLL, so you will have to manually generate it in simulation.
    always_ff @ (posedge VGA_CLK)
    begin
        if (Reset)
        begin
            VGA_HS <= 1'b0;
            VGA_VS <= 1'b0;
            VGA_BLANK_N <= 1'b0;
            h_counter <= 10'd0;
            v_counter <= 10'd0;
        end
        else
        begin
            VGA_HS <= VGA_HS_in;
            VGA_VS <= VGA_VS_in;
            VGA_BLANK_N <= VGA_BLANK_N_in;
            h_counter <= h_counter_in;
            v_counter <= v_counter_in;
        end
    end
    
    always_comb
    begin
        // horizontal and vertical counter
        h_counter_in = h_counter + 10'd1;
        v_counter_in = v_counter;
        if(h_counter + 10'd1 == H_TOTAL)
        begin
            h_counter_in = 10'd0;
            if(v_counter + 10'd1 == V_TOTAL)
                v_counter_in = 10'd0;
            else
                v_counter_in = v_counter + 10'd1;
        end
        // Horizontal sync pulse is 96 pixels long at pixels 656-752
        // (Signal is registered to ensure clean output waveform)
        VGA_HS_in = 1'b1;
        if(h_counter_in >= 10'd656 && h_counter_in < 10'd752)
            VGA_HS_in = 1'b0;
        // Vertical sync pulse is 2 lines (800 pixels each) long at line 490-491
        //(Signal is registered to ensure clean output waveform)
        VGA_VS_in = 1'b1;
        if(v_counter_in >= 10'd490 && v_counter_in < 10'd492)
            VGA_VS_in = 1'b0;
        // Display pixels (inhibit blanking) between horizontal 0-639 and vertical 0-479 (640x480)
        VGA_BLANK_N_in = 1'b0;
        if(h_counter_in < 10'd640 && v_counter_in < 10'd480)
            VGA_BLANK_N_in = 1'b1;
    end
    
endmodule


module VGA_mapper(
    input logic CLK, RESET,
    input logic [11:0] VGA_ADDR,
    input logic [7:0] VGA_WRITEDATA,
    output logic [7:0] VGA_READDATA,
    input logic VGA_WRITE, VGA_CS, VGA_BYTE_EN, VGA_READ,
    input logic VGA_BLANK_N,
    output logic [7:0] VGA_R, VGA_G, VGA_B
);

    logic [7:0] ram1_data, ram2_data;
    logic ram1_we, ram2_we;
    logic current_ram = 0;
    logic needs_write = 0;
    logic needs_write_next;

    logic [10:0] draw_counter = 0;
    logic [1:0] rgb_counter = 0;

    logic [7:0] signal_reg, signal_reg_next;

    vga_ram #(0) ram1(.output_data(ram1_data),
        .input_data(VGA_WRITEDATA), 
        .write_address(VGA_ADDR[10:0]), .read_address(draw_counter),
        .we(ram1_we), .clk(CLK));

    vga_ram #(1) ram2(.output_data(ram2_data),
        .input_data(VGA_WRITEDATA), 
        .write_address(VGA_ADDR[10:0]), .read_address(draw_counter),
        .we(ram2_we), .clk(CLK));


    always_comb begin

        if(VGA_ADDR == 1920) begin
            ram1_we = 1'b0;
            ram2_we = 1'b0;
            needs_write_next = needs_write;
        end else if (VGA_ADDR == 1921) begin
            ram1_we = 1'b0;
            ram2_we = 1'b0;
            if(VGA_CS & VGA_WRITE & VGA_BYTE_EN)
                needs_write_next = 0;
            else
                needs_write_next = needs_write;
        end else if(VGA_ADDR[11] == 0) begin
            ram1_we = VGA_WRITE & VGA_CS & VGA_BYTE_EN;
            ram2_we = 1'b0;
            needs_write_next = needs_write;
        end else if(VGA_ADDR[11] == 1) begin
            ram2_we = VGA_WRITE & VGA_CS & VGA_BYTE_EN;
            ram1_we = 1'b0;
            needs_write_next = needs_write;
        end else begin
            ram1_we = 1'b0;
            ram2_we = 1'b0;
            needs_write_next = needs_write;
        end

        if(draw_counter == 1919)
            needs_write_next = 1;
        else
            needs_write_next = needs_write;
        
        if(VGA_READ & VGA_CS) begin
            if(VGA_ADDR == 1920) 
                VGA_READDATA = {7'b0000000, current_ram};
            else if (VGA_ADDR == 1921)
                VGA_READDATA = {7'b0000000, needs_write};
            else
                VGA_READDATA = 8'bzzzzzzzz;
        end else
            VGA_READDATA = 8'bzzzzzzzz;


    end

     always_ff @(posedge CLK) begin

         if (RESET)
             needs_write <= 0;
         else
             needs_write <= needs_write_next;

         if (RESET)
             draw_counter <= 0;
         else if(draw_counter == 1919) begin
             draw_counter <= 0;
             if(current_ram == 0)
                 current_ram <= 1;
             else
                 current_ram <= 0;
         end
         else if(VGA_BLANK_N)
             draw_counter <= (draw_counter+1);
         else
             draw_counter <= draw_counter;
 
         if (RESET || (VGA_BLANK_N == 0))
             rgb_counter <= 0;
         else if(rgb_counter == 2)
             rgb_counter <= 0;
         else if(VGA_BLANK_N)
             rgb_counter <= (rgb_counter + 1);
         else
             rgb_counter <= rgb_counter;
 
         if(current_ram == 0) begin
             if(rgb_counter == 0)
                 VGA_R <= ram1_data;
             else if (rgb_counter == 1)
                 VGA_G <= ram1_data;
             else
                 VGA_B <= ram1_data;
         end else begin
             if(rgb_counter == 0)
                 VGA_R <= ram2_data;
             else if (rgb_counter == 1)
                 VGA_G <= ram2_data;
             else
                 VGA_B <= ram2_data;
         end
 
 
     end
     
 
endmodule

module vga_ram #(parameter ram_num = 0)(
    output logic [7:0] output_data,
    input logic [7:0] input_data,
    input [10:0] write_address, read_address,
    input we, clk
);

logic [7:0] mem[1920];

initial
begin
    if(ram_num == 0) begin
        $display("Reading ram 0");
        $readmemh("vga_ram0.txt", mem);
    end else if(ram_num == 1) begin
        $display("Reading ram 1");
        $readmemh("vga_ram1.txt", mem);
    end else begin
        $display("Unknown ram number----------------------");
    end
end

always_ff @ (posedge clk) begin
    if (we)
        mem[write_address] <= input_data;
    output_data <= mem[read_address];

end
endmodule
