// final_soc.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module final_soc (
		input  wire        clk_clk,                //             clk.clk
		output wire [7:0]  keycode_export,         //         keycode.export
		output wire [1:0]  otg_hpi_address_export, // otg_hpi_address.export
		output wire        otg_hpi_cs_export,      //      otg_hpi_cs.export
		input  wire [15:0] otg_hpi_data_in_port,   //    otg_hpi_data.in_port
		output wire [15:0] otg_hpi_data_out_port,  //                .out_port
		output wire        otg_hpi_r_export,       //       otg_hpi_r.export
		output wire        otg_hpi_reset_export,   //   otg_hpi_reset.export
		output wire        otg_hpi_w_export,       //       otg_hpi_w.export
		input  wire        reset_reset_n,          //           reset.reset_n
		output wire        sdram_clk_clk,          //       sdram_clk.clk
		output wire [12:0] sdram_wire_addr,        //      sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,          //                .ba
		output wire        sdram_wire_cas_n,       //                .cas_n
		output wire        sdram_wire_cke,         //                .cke
		output wire        sdram_wire_cs_n,        //                .cs_n
		inout  wire [31:0] sdram_wire_dq,          //                .dq
		output wire [3:0]  sdram_wire_dqm,         //                .dqm
		output wire        sdram_wire_ras_n,       //                .ras_n
		output wire        sdram_wire_we_n,        //                .we_n
		output wire        vga_CLK,                //             vga.CLK
		output wire        vga_HS,                 //                .HS
		output wire        vga_VS,                 //                .VS
		output wire        vga_BLANK,              //                .BLANK
		output wire        vga_SYNC,               //                .SYNC
		output wire [7:0]  vga_R,                  //                .R
		output wire [7:0]  vga_G,                  //                .G
		output wire [7:0]  vga_B                   //                .B
	);

	wire         pixel_out_buffer_avalon_dc_buffer_source_valid;              // pixel_out_buffer:stream_out_valid -> vga_resampler:stream_in_valid
	wire  [31:0] pixel_out_buffer_avalon_dc_buffer_source_data;               // pixel_out_buffer:stream_out_data -> vga_resampler:stream_in_data
	wire         pixel_out_buffer_avalon_dc_buffer_source_ready;              // vga_resampler:stream_in_ready -> pixel_out_buffer:stream_out_ready
	wire         pixel_out_buffer_avalon_dc_buffer_source_startofpacket;      // pixel_out_buffer:stream_out_startofpacket -> vga_resampler:stream_in_startofpacket
	wire         pixel_out_buffer_avalon_dc_buffer_source_endofpacket;        // pixel_out_buffer:stream_out_endofpacket -> vga_resampler:stream_in_endofpacket
	wire         pixel_dma_avalon_pixel_source_valid;                         // pixel_dma:stream_valid -> pixel_out_buffer:stream_in_valid
	wire  [31:0] pixel_dma_avalon_pixel_source_data;                          // pixel_dma:stream_data -> pixel_out_buffer:stream_in_data
	wire         pixel_dma_avalon_pixel_source_ready;                         // pixel_out_buffer:stream_in_ready -> pixel_dma:stream_ready
	wire         pixel_dma_avalon_pixel_source_startofpacket;                 // pixel_dma:stream_startofpacket -> pixel_out_buffer:stream_in_startofpacket
	wire         pixel_dma_avalon_pixel_source_endofpacket;                   // pixel_dma:stream_endofpacket -> pixel_out_buffer:stream_in_endofpacket
	wire         vga_resampler_avalon_rgb_source_valid;                       // vga_resampler:stream_out_valid -> vga_scaler:stream_in_valid
	wire  [29:0] vga_resampler_avalon_rgb_source_data;                        // vga_resampler:stream_out_data -> vga_scaler:stream_in_data
	wire         vga_resampler_avalon_rgb_source_ready;                       // vga_scaler:stream_in_ready -> vga_resampler:stream_out_ready
	wire         vga_resampler_avalon_rgb_source_startofpacket;               // vga_resampler:stream_out_startofpacket -> vga_scaler:stream_in_startofpacket
	wire         vga_resampler_avalon_rgb_source_endofpacket;                 // vga_resampler:stream_out_endofpacket -> vga_scaler:stream_in_endofpacket
	wire         pll_c0_clk;                                                  // PLL:c0 -> [SDRAM:clk, mm_interconnect_0:PLL_c0_clk, rst_controller_001:clk]
	wire         pll_c2_clk;                                                  // PLL:c2 -> [avalon_st_adapter:in_clk_0_clk, mm_interconnect_0:PLL_c2_clk, pixel_out_buffer:clk_stream_out, rst_controller_002:clk, vga_controller:clk, vga_resampler:clk, vga_scaler:clk]
	wire         gpu_core_0_gpu_master_chipselect;                            // GPU_CORE_0:GPU_MASTER_chipselect -> mm_interconnect_0:GPU_CORE_0_GPU_MASTER_chipselect
	wire  [31:0] gpu_core_0_gpu_master_readdata;                              // mm_interconnect_0:GPU_CORE_0_GPU_MASTER_readdata -> GPU_CORE_0:GPU_MASTER_readdata
	wire         gpu_core_0_gpu_master_waitrequest;                           // mm_interconnect_0:GPU_CORE_0_GPU_MASTER_waitrequest -> GPU_CORE_0:GPU_MASTER_waitrequest
	wire  [31:0] gpu_core_0_gpu_master_address;                               // GPU_CORE_0:GPU_MASTER_address -> mm_interconnect_0:GPU_CORE_0_GPU_MASTER_address
	wire         gpu_core_0_gpu_master_read;                                  // GPU_CORE_0:GPU_MASTER_read -> mm_interconnect_0:GPU_CORE_0_GPU_MASTER_read
	wire         gpu_core_0_gpu_master_readdatavalid;                         // mm_interconnect_0:GPU_CORE_0_GPU_MASTER_readdatavalid -> GPU_CORE_0:GPU_MASTER_readdatavalid
	wire   [1:0] gpu_core_0_gpu_master_response;                              // mm_interconnect_0:GPU_CORE_0_GPU_MASTER_response -> GPU_CORE_0:GPU_MASTER_response
	wire         gpu_core_0_gpu_master_write;                                 // GPU_CORE_0:GPU_MASTER_write -> mm_interconnect_0:GPU_CORE_0_GPU_MASTER_write
	wire  [31:0] gpu_core_0_gpu_master_writedata;                             // GPU_CORE_0:GPU_MASTER_writedata -> mm_interconnect_0:GPU_CORE_0_GPU_MASTER_writedata
	wire         gpu_core_0_gpu_master_writeresponsevalid;                    // mm_interconnect_0:GPU_CORE_0_GPU_MASTER_writeresponsevalid -> GPU_CORE_0:GPU_MASTER_writeresponsevalid
	wire  [31:0] nios2_data_master_readdata;                                  // mm_interconnect_0:NIOS2_data_master_readdata -> NIOS2:d_readdata
	wire         nios2_data_master_waitrequest;                               // mm_interconnect_0:NIOS2_data_master_waitrequest -> NIOS2:d_waitrequest
	wire         nios2_data_master_debugaccess;                               // NIOS2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS2_data_master_debugaccess
	wire  [27:0] nios2_data_master_address;                                   // NIOS2:d_address -> mm_interconnect_0:NIOS2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                                // NIOS2:d_byteenable -> mm_interconnect_0:NIOS2_data_master_byteenable
	wire         nios2_data_master_read;                                      // NIOS2:d_read -> mm_interconnect_0:NIOS2_data_master_read
	wire         nios2_data_master_write;                                     // NIOS2:d_write -> mm_interconnect_0:NIOS2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                                 // NIOS2:d_writedata -> mm_interconnect_0:NIOS2_data_master_writedata
	wire         pixel_dma_avalon_pixel_dma_master_waitrequest;               // mm_interconnect_0:pixel_dma_avalon_pixel_dma_master_waitrequest -> pixel_dma:master_waitrequest
	wire  [31:0] pixel_dma_avalon_pixel_dma_master_readdata;                  // mm_interconnect_0:pixel_dma_avalon_pixel_dma_master_readdata -> pixel_dma:master_readdata
	wire  [31:0] pixel_dma_avalon_pixel_dma_master_address;                   // pixel_dma:master_address -> mm_interconnect_0:pixel_dma_avalon_pixel_dma_master_address
	wire         pixel_dma_avalon_pixel_dma_master_read;                      // pixel_dma:master_read -> mm_interconnect_0:pixel_dma_avalon_pixel_dma_master_read
	wire         pixel_dma_avalon_pixel_dma_master_readdatavalid;             // mm_interconnect_0:pixel_dma_avalon_pixel_dma_master_readdatavalid -> pixel_dma:master_readdatavalid
	wire         pixel_dma_avalon_pixel_dma_master_lock;                      // pixel_dma:master_arbiterlock -> mm_interconnect_0:pixel_dma_avalon_pixel_dma_master_lock
	wire  [31:0] nios2_instruction_master_readdata;                           // mm_interconnect_0:NIOS2_instruction_master_readdata -> NIOS2:i_readdata
	wire         nios2_instruction_master_waitrequest;                        // mm_interconnect_0:NIOS2_instruction_master_waitrequest -> NIOS2:i_waitrequest
	wire  [27:0] nios2_instruction_master_address;                            // NIOS2:i_address -> mm_interconnect_0:NIOS2_instruction_master_address
	wire         nios2_instruction_master_read;                               // NIOS2:i_read -> mm_interconnect_0:NIOS2_instruction_master_read
	wire         mm_interconnect_0_frame_buffer_s1_chipselect;                // mm_interconnect_0:frame_buffer_s1_chipselect -> frame_buffer:chipselect
	wire  [31:0] mm_interconnect_0_frame_buffer_s1_readdata;                  // frame_buffer:readdata -> mm_interconnect_0:frame_buffer_s1_readdata
	wire  [16:0] mm_interconnect_0_frame_buffer_s1_address;                   // mm_interconnect_0:frame_buffer_s1_address -> frame_buffer:address
	wire   [3:0] mm_interconnect_0_frame_buffer_s1_byteenable;                // mm_interconnect_0:frame_buffer_s1_byteenable -> frame_buffer:byteenable
	wire         mm_interconnect_0_frame_buffer_s1_write;                     // mm_interconnect_0:frame_buffer_s1_write -> frame_buffer:write
	wire  [31:0] mm_interconnect_0_frame_buffer_s1_writedata;                 // mm_interconnect_0:frame_buffer_s1_writedata -> frame_buffer:writedata
	wire         mm_interconnect_0_frame_buffer_s1_clken;                     // mm_interconnect_0:frame_buffer_s1_clken -> frame_buffer:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                       // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                         // SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                      // SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                          // mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                             // mm_interconnect_0:SDRAM_s1_read -> SDRAM:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                       // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                    // SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                            // mm_interconnect_0:SDRAM_s1_write -> SDRAM:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                        // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	wire         mm_interconnect_0_gpu_core_0_gpu_slave_chipselect;           // mm_interconnect_0:GPU_CORE_0_GPU_SLAVE_chipselect -> GPU_CORE_0:GPU_SLAVE_chipselect
	wire  [31:0] mm_interconnect_0_gpu_core_0_gpu_slave_readdata;             // GPU_CORE_0:GPU_SLAVE_readdata -> mm_interconnect_0:GPU_CORE_0_GPU_SLAVE_readdata
	wire  [10:0] mm_interconnect_0_gpu_core_0_gpu_slave_address;              // mm_interconnect_0:GPU_CORE_0_GPU_SLAVE_address -> GPU_CORE_0:GPU_SLAVE_address
	wire         mm_interconnect_0_gpu_core_0_gpu_slave_read;                 // mm_interconnect_0:GPU_CORE_0_GPU_SLAVE_read -> GPU_CORE_0:GPU_SLAVE_read
	wire         mm_interconnect_0_gpu_core_0_gpu_slave_write;                // mm_interconnect_0:GPU_CORE_0_GPU_SLAVE_write -> GPU_CORE_0:GPU_SLAVE_write
	wire  [31:0] mm_interconnect_0_gpu_core_0_gpu_slave_writedata;            // mm_interconnect_0:GPU_CORE_0_GPU_SLAVE_writedata -> GPU_CORE_0:GPU_SLAVE_writedata
	wire  [31:0] mm_interconnect_0_pixel_dma_avalon_control_slave_readdata;   // pixel_dma:slave_readdata -> mm_interconnect_0:pixel_dma_avalon_control_slave_readdata
	wire   [1:0] mm_interconnect_0_pixel_dma_avalon_control_slave_address;    // mm_interconnect_0:pixel_dma_avalon_control_slave_address -> pixel_dma:slave_address
	wire         mm_interconnect_0_pixel_dma_avalon_control_slave_read;       // mm_interconnect_0:pixel_dma_avalon_control_slave_read -> pixel_dma:slave_read
	wire   [3:0] mm_interconnect_0_pixel_dma_avalon_control_slave_byteenable; // mm_interconnect_0:pixel_dma_avalon_control_slave_byteenable -> pixel_dma:slave_byteenable
	wire         mm_interconnect_0_pixel_dma_avalon_control_slave_write;      // mm_interconnect_0:pixel_dma_avalon_control_slave_write -> pixel_dma:slave_write
	wire  [31:0] mm_interconnect_0_pixel_dma_avalon_control_slave_writedata;  // mm_interconnect_0:pixel_dma_avalon_control_slave_writedata -> pixel_dma:slave_writedata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_vga_resampler_avalon_rgb_slave_readdata;   // vga_resampler:slave_readdata -> mm_interconnect_0:vga_resampler_avalon_rgb_slave_readdata
	wire         mm_interconnect_0_vga_resampler_avalon_rgb_slave_read;       // mm_interconnect_0:vga_resampler_avalon_rgb_slave_read -> vga_resampler:slave_read
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;            // NIOS2:debug_mem_slave_readdata -> mm_interconnect_0:NIOS2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;         // NIOS2:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;         // mm_interconnect_0:NIOS2_debug_mem_slave_debugaccess -> NIOS2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;             // mm_interconnect_0:NIOS2_debug_mem_slave_address -> NIOS2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;                // mm_interconnect_0:NIOS2_debug_mem_slave_read -> NIOS2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;          // mm_interconnect_0:NIOS2_debug_mem_slave_byteenable -> NIOS2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;               // mm_interconnect_0:NIOS2_debug_mem_slave_write -> NIOS2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;           // mm_interconnect_0:NIOS2_debug_mem_slave_writedata -> NIOS2:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_pll_pll_slave_readdata;                    // PLL:readdata -> mm_interconnect_0:PLL_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_pll_pll_slave_address;                     // mm_interconnect_0:PLL_pll_slave_address -> PLL:address
	wire         mm_interconnect_0_pll_pll_slave_read;                        // mm_interconnect_0:PLL_pll_slave_read -> PLL:read
	wire         mm_interconnect_0_pll_pll_slave_write;                       // mm_interconnect_0:PLL_pll_slave_write -> PLL:write
	wire  [31:0] mm_interconnect_0_pll_pll_slave_writedata;                   // mm_interconnect_0:PLL_pll_slave_writedata -> PLL:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_keycode_s1_chipselect;                     // mm_interconnect_0:keycode_s1_chipselect -> keycode:chipselect
	wire  [31:0] mm_interconnect_0_keycode_s1_readdata;                       // keycode:readdata -> mm_interconnect_0:keycode_s1_readdata
	wire   [1:0] mm_interconnect_0_keycode_s1_address;                        // mm_interconnect_0:keycode_s1_address -> keycode:address
	wire         mm_interconnect_0_keycode_s1_write;                          // mm_interconnect_0:keycode_s1_write -> keycode:write_n
	wire  [31:0] mm_interconnect_0_keycode_s1_writedata;                      // mm_interconnect_0:keycode_s1_writedata -> keycode:writedata
	wire         mm_interconnect_0_otg_hpi_address_s1_chipselect;             // mm_interconnect_0:otg_hpi_address_s1_chipselect -> otg_hpi_address:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_address_s1_readdata;               // otg_hpi_address:readdata -> mm_interconnect_0:otg_hpi_address_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_address_s1_address;                // mm_interconnect_0:otg_hpi_address_s1_address -> otg_hpi_address:address
	wire         mm_interconnect_0_otg_hpi_address_s1_write;                  // mm_interconnect_0:otg_hpi_address_s1_write -> otg_hpi_address:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_address_s1_writedata;              // mm_interconnect_0:otg_hpi_address_s1_writedata -> otg_hpi_address:writedata
	wire         mm_interconnect_0_otg_hpi_data_s1_chipselect;                // mm_interconnect_0:otg_hpi_data_s1_chipselect -> otg_hpi_data:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_data_s1_readdata;                  // otg_hpi_data:readdata -> mm_interconnect_0:otg_hpi_data_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_data_s1_address;                   // mm_interconnect_0:otg_hpi_data_s1_address -> otg_hpi_data:address
	wire         mm_interconnect_0_otg_hpi_data_s1_write;                     // mm_interconnect_0:otg_hpi_data_s1_write -> otg_hpi_data:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_data_s1_writedata;                 // mm_interconnect_0:otg_hpi_data_s1_writedata -> otg_hpi_data:writedata
	wire         mm_interconnect_0_otg_hpi_r_s1_chipselect;                   // mm_interconnect_0:otg_hpi_r_s1_chipselect -> otg_hpi_r:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_r_s1_readdata;                     // otg_hpi_r:readdata -> mm_interconnect_0:otg_hpi_r_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_r_s1_address;                      // mm_interconnect_0:otg_hpi_r_s1_address -> otg_hpi_r:address
	wire         mm_interconnect_0_otg_hpi_r_s1_write;                        // mm_interconnect_0:otg_hpi_r_s1_write -> otg_hpi_r:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_r_s1_writedata;                    // mm_interconnect_0:otg_hpi_r_s1_writedata -> otg_hpi_r:writedata
	wire         mm_interconnect_0_otg_hpi_w_s1_chipselect;                   // mm_interconnect_0:otg_hpi_w_s1_chipselect -> otg_hpi_w:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_w_s1_readdata;                     // otg_hpi_w:readdata -> mm_interconnect_0:otg_hpi_w_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_w_s1_address;                      // mm_interconnect_0:otg_hpi_w_s1_address -> otg_hpi_w:address
	wire         mm_interconnect_0_otg_hpi_w_s1_write;                        // mm_interconnect_0:otg_hpi_w_s1_write -> otg_hpi_w:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_w_s1_writedata;                    // mm_interconnect_0:otg_hpi_w_s1_writedata -> otg_hpi_w:writedata
	wire         mm_interconnect_0_otg_hpi_cs_s1_chipselect;                  // mm_interconnect_0:otg_hpi_cs_s1_chipselect -> otg_hpi_cs:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_cs_s1_readdata;                    // otg_hpi_cs:readdata -> mm_interconnect_0:otg_hpi_cs_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_cs_s1_address;                     // mm_interconnect_0:otg_hpi_cs_s1_address -> otg_hpi_cs:address
	wire         mm_interconnect_0_otg_hpi_cs_s1_write;                       // mm_interconnect_0:otg_hpi_cs_s1_write -> otg_hpi_cs:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_cs_s1_writedata;                   // mm_interconnect_0:otg_hpi_cs_s1_writedata -> otg_hpi_cs:writedata
	wire         mm_interconnect_0_otg_hpi_reset_s1_chipselect;               // mm_interconnect_0:otg_hpi_reset_s1_chipselect -> otg_hpi_reset:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_reset_s1_readdata;                 // otg_hpi_reset:readdata -> mm_interconnect_0:otg_hpi_reset_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_reset_s1_address;                  // mm_interconnect_0:otg_hpi_reset_s1_address -> otg_hpi_reset:address
	wire         mm_interconnect_0_otg_hpi_reset_s1_write;                    // mm_interconnect_0:otg_hpi_reset_s1_write -> otg_hpi_reset:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_reset_s1_writedata;                // mm_interconnect_0:otg_hpi_reset_s1_writedata -> otg_hpi_reset:writedata
	wire         mm_interconnect_0_frame_buffer_s2_chipselect;                // mm_interconnect_0:frame_buffer_s2_chipselect -> frame_buffer:chipselect2
	wire  [31:0] mm_interconnect_0_frame_buffer_s2_readdata;                  // frame_buffer:readdata2 -> mm_interconnect_0:frame_buffer_s2_readdata
	wire  [16:0] mm_interconnect_0_frame_buffer_s2_address;                   // mm_interconnect_0:frame_buffer_s2_address -> frame_buffer:address2
	wire   [3:0] mm_interconnect_0_frame_buffer_s2_byteenable;                // mm_interconnect_0:frame_buffer_s2_byteenable -> frame_buffer:byteenable2
	wire         mm_interconnect_0_frame_buffer_s2_write;                     // mm_interconnect_0:frame_buffer_s2_write -> frame_buffer:write2
	wire  [31:0] mm_interconnect_0_frame_buffer_s2_writedata;                 // mm_interconnect_0:frame_buffer_s2_writedata -> frame_buffer:writedata2
	wire         mm_interconnect_0_frame_buffer_s2_clken;                     // mm_interconnect_0:frame_buffer_s2_clken -> frame_buffer:clken2
	wire         irq_mapper_receiver0_irq;                                    // timer_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_irq_irq;                                               // irq_mapper:sender_irq -> NIOS2:irq
	wire         vga_scaler_avalon_scaler_source_valid;                       // vga_scaler:stream_out_valid -> avalon_st_adapter:in_0_valid
	wire  [29:0] vga_scaler_avalon_scaler_source_data;                        // vga_scaler:stream_out_data -> avalon_st_adapter:in_0_data
	wire         vga_scaler_avalon_scaler_source_ready;                       // avalon_st_adapter:in_0_ready -> vga_scaler:stream_out_ready
	wire   [1:0] vga_scaler_avalon_scaler_source_channel;                     // vga_scaler:stream_out_channel -> avalon_st_adapter:in_0_channel
	wire         vga_scaler_avalon_scaler_source_startofpacket;               // vga_scaler:stream_out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire         vga_scaler_avalon_scaler_source_endofpacket;                 // vga_scaler:stream_out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire         avalon_st_adapter_out_0_valid;                               // avalon_st_adapter:out_0_valid -> vga_controller:valid
	wire  [29:0] avalon_st_adapter_out_0_data;                                // avalon_st_adapter:out_0_data -> vga_controller:data
	wire         avalon_st_adapter_out_0_ready;                               // vga_controller:ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                       // avalon_st_adapter:out_0_startofpacket -> vga_controller:startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                         // avalon_st_adapter:out_0_endofpacket -> vga_controller:endofpacket
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [GPU_CORE_0:RESET_reset, NIOS2:reset_n, PLL:reset, frame_buffer:reset, frame_buffer:reset2, irq_mapper:reset, jtag_uart_0:rst_n, keycode:reset_n, mm_interconnect_0:GPU_CORE_0_RESET_reset_bridge_in_reset_reset, otg_hpi_address:reset_n, otg_hpi_cs:reset_n, otg_hpi_data:reset_n, otg_hpi_r:reset_n, otg_hpi_reset:reset_n, otg_hpi_w:reset_n, pixel_dma:reset, pixel_out_buffer:reset_stream_in, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [NIOS2:reset_req, frame_buffer:reset_req, frame_buffer:reset_req2, rst_translator:reset_req_in]
	wire         nios2_debug_reset_request_reset;                             // NIOS2:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [SDRAM:reset_n, mm_interconnect_0:SDRAM_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;                          // rst_controller_002:reset_out -> [avalon_st_adapter:in_rst_0_reset, mm_interconnect_0:vga_resampler_reset_reset_bridge_in_reset_reset, pixel_out_buffer:reset_stream_out, vga_controller:reset, vga_resampler:reset, vga_scaler:reset]
	wire         rst_controller_003_reset_out_reset;                          // rst_controller_003:reset_out -> [mm_interconnect_0:timer_0_reset_reset_bridge_in_reset_reset, timer_0:reset_n]

	avalon_gpu_interface gpu_core_0 (
		.CLK_clk                       (clk_clk),                                           //        CLK.clk
		.RESET_reset                   (rst_controller_reset_out_reset),                    //      RESET.reset
		.GPU_SLAVE_read                (mm_interconnect_0_gpu_core_0_gpu_slave_read),       //  GPU_SLAVE.read
		.GPU_SLAVE_readdata            (mm_interconnect_0_gpu_core_0_gpu_slave_readdata),   //           .readdata
		.GPU_SLAVE_write               (mm_interconnect_0_gpu_core_0_gpu_slave_write),      //           .write
		.GPU_SLAVE_writedata           (mm_interconnect_0_gpu_core_0_gpu_slave_writedata),  //           .writedata
		.GPU_SLAVE_address             (mm_interconnect_0_gpu_core_0_gpu_slave_address),    //           .address
		.GPU_SLAVE_chipselect          (mm_interconnect_0_gpu_core_0_gpu_slave_chipselect), //           .chipselect
		.GPU_MASTER_address            (gpu_core_0_gpu_master_address),                     // GPU_MASTER.address
		.GPU_MASTER_read               (gpu_core_0_gpu_master_read),                        //           .read
		.GPU_MASTER_readdata           (gpu_core_0_gpu_master_readdata),                    //           .readdata
		.GPU_MASTER_chipselect         (gpu_core_0_gpu_master_chipselect),                  //           .chipselect
		.GPU_MASTER_readdatavalid      (gpu_core_0_gpu_master_readdatavalid),               //           .readdatavalid
		.GPU_MASTER_writeresponsevalid (gpu_core_0_gpu_master_writeresponsevalid),          //           .writeresponsevalid
		.GPU_MASTER_write              (gpu_core_0_gpu_master_write),                       //           .write
		.GPU_MASTER_writedata          (gpu_core_0_gpu_master_writedata),                   //           .writedata
		.GPU_MASTER_response           (gpu_core_0_gpu_master_response),                    //           .response
		.GPU_MASTER_waitrequest        (gpu_core_0_gpu_master_waitrequest)                  //           .waitrequest
	);

	final_soc_NIOS2 nios2 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	final_soc_PLL pll (
		.clk                (clk_clk),                                   //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),            // inclk_interface_reset.reset
		.read               (mm_interconnect_0_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_pll_pll_slave_writedata), //                      .writedata
		.c0                 (pll_c0_clk),                                //                    c0.clk
		.c1                 (sdram_clk_clk),                             //                    c1.clk
		.c2                 (pll_c2_clk),                                //                    c2.clk
		.c3                 (),                                          //                    c3.clk
		.c4                 (),                                          //                    c4.clk
		.scandone           (),                                          //           (terminated)
		.scandataout        (),                                          //           (terminated)
		.areset             (1'b0),                                      //           (terminated)
		.locked             (),                                          //           (terminated)
		.phasedone          (),                                          //           (terminated)
		.phasecounterselect (4'b0000),                                   //           (terminated)
		.phaseupdown        (1'b0),                                      //           (terminated)
		.phasestep          (1'b0),                                      //           (terminated)
		.scanclk            (1'b0),                                      //           (terminated)
		.scanclkena         (1'b0),                                      //           (terminated)
		.scandata           (1'b0),                                      //           (terminated)
		.configupdate       (1'b0)                                       //           (terminated)
	);

	final_soc_SDRAM sdram (
		.clk            (pll_c0_clk),                               //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	final_soc_frame_buffer frame_buffer (
		.clk         (clk_clk),                                      //   clk1.clk
		.address     (mm_interconnect_0_frame_buffer_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_frame_buffer_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_frame_buffer_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_frame_buffer_s1_write),      //       .write
		.readdata    (mm_interconnect_0_frame_buffer_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_frame_buffer_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_frame_buffer_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),               // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),           //       .reset_req
		.address2    (mm_interconnect_0_frame_buffer_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_frame_buffer_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_frame_buffer_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_frame_buffer_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_frame_buffer_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_frame_buffer_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_frame_buffer_s2_byteenable), //       .byteenable
		.clk2        (clk_clk),                                      //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),               // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req),           //       .reset_req
		.freeze      (1'b0)                                          // (terminated)
	);

	final_soc_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	final_soc_keycode keycode (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_keycode_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keycode_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keycode_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keycode_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keycode_s1_readdata),   //                    .readdata
		.out_port   (keycode_export)                           // external_connection.export
	);

	final_soc_otg_hpi_address otg_hpi_address (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_address_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_address_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_address_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_address_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_address_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_address_export)                           // external_connection.export
	);

	final_soc_otg_hpi_cs otg_hpi_cs (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_cs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_cs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_cs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_cs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_cs_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_cs_export)                           // external_connection.export
	);

	final_soc_otg_hpi_data otg_hpi_data (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_data_s1_readdata),   //                    .readdata
		.in_port    (otg_hpi_data_in_port),                         // external_connection.export
		.out_port   (otg_hpi_data_out_port)                         //                    .export
	);

	final_soc_otg_hpi_cs otg_hpi_r (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_r_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_r_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_r_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_r_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_r_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_r_export)                           // external_connection.export
	);

	final_soc_otg_hpi_cs otg_hpi_reset (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_reset_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_reset_export)                           // external_connection.export
	);

	final_soc_otg_hpi_cs otg_hpi_w (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_w_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_w_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_w_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_w_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_w_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_w_export)                           // external_connection.export
	);

	final_soc_pixel_dma pixel_dma (
		.clk                  (clk_clk),                                                     //                     clk.clk
		.reset                (rst_controller_reset_out_reset),                              //                   reset.reset
		.master_readdatavalid (pixel_dma_avalon_pixel_dma_master_readdatavalid),             // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (pixel_dma_avalon_pixel_dma_master_waitrequest),               //                        .waitrequest
		.master_address       (pixel_dma_avalon_pixel_dma_master_address),                   //                        .address
		.master_arbiterlock   (pixel_dma_avalon_pixel_dma_master_lock),                      //                        .lock
		.master_read          (pixel_dma_avalon_pixel_dma_master_read),                      //                        .read
		.master_readdata      (pixel_dma_avalon_pixel_dma_master_readdata),                  //                        .readdata
		.slave_address        (mm_interconnect_0_pixel_dma_avalon_control_slave_address),    //    avalon_control_slave.address
		.slave_byteenable     (mm_interconnect_0_pixel_dma_avalon_control_slave_byteenable), //                        .byteenable
		.slave_read           (mm_interconnect_0_pixel_dma_avalon_control_slave_read),       //                        .read
		.slave_write          (mm_interconnect_0_pixel_dma_avalon_control_slave_write),      //                        .write
		.slave_writedata      (mm_interconnect_0_pixel_dma_avalon_control_slave_writedata),  //                        .writedata
		.slave_readdata       (mm_interconnect_0_pixel_dma_avalon_control_slave_readdata),   //                        .readdata
		.stream_ready         (pixel_dma_avalon_pixel_source_ready),                         //     avalon_pixel_source.ready
		.stream_startofpacket (pixel_dma_avalon_pixel_source_startofpacket),                 //                        .startofpacket
		.stream_endofpacket   (pixel_dma_avalon_pixel_source_endofpacket),                   //                        .endofpacket
		.stream_valid         (pixel_dma_avalon_pixel_source_valid),                         //                        .valid
		.stream_data          (pixel_dma_avalon_pixel_source_data)                           //                        .data
	);

	final_soc_pixel_out_buffer pixel_out_buffer (
		.clk_stream_in            (clk_clk),                                                //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_reset_out_reset),                         //         reset_stream_in.reset
		.clk_stream_out           (pll_c2_clk),                                             //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_002_reset_out_reset),                     //        reset_stream_out.reset
		.stream_in_ready          (pixel_dma_avalon_pixel_source_ready),                    //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (pixel_dma_avalon_pixel_source_startofpacket),            //                        .startofpacket
		.stream_in_endofpacket    (pixel_dma_avalon_pixel_source_endofpacket),              //                        .endofpacket
		.stream_in_valid          (pixel_dma_avalon_pixel_source_valid),                    //                        .valid
		.stream_in_data           (pixel_dma_avalon_pixel_source_data),                     //                        .data
		.stream_out_ready         (pixel_out_buffer_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (pixel_out_buffer_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (pixel_out_buffer_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (pixel_out_buffer_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (pixel_out_buffer_avalon_dc_buffer_source_data)           //                        .data
	);

	final_soc_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                 //   irq.irq
	);

	final_soc_vga_controller vga_controller (
		.clk           (pll_c2_clk),                            //                clk.clk
		.reset         (rst_controller_002_reset_out_reset),    //              reset.reset
		.data          (avalon_st_adapter_out_0_data),          //    avalon_vga_sink.data
		.startofpacket (avalon_st_adapter_out_0_startofpacket), //                   .startofpacket
		.endofpacket   (avalon_st_adapter_out_0_endofpacket),   //                   .endofpacket
		.valid         (avalon_st_adapter_out_0_valid),         //                   .valid
		.ready         (avalon_st_adapter_out_0_ready),         //                   .ready
		.VGA_CLK       (vga_CLK),                               // external_interface.export
		.VGA_HS        (vga_HS),                                //                   .export
		.VGA_VS        (vga_VS),                                //                   .export
		.VGA_BLANK     (vga_BLANK),                             //                   .export
		.VGA_SYNC      (vga_SYNC),                              //                   .export
		.VGA_R         (vga_R),                                 //                   .export
		.VGA_G         (vga_G),                                 //                   .export
		.VGA_B         (vga_B)                                  //                   .export
	);

	final_soc_vga_resampler vga_resampler (
		.clk                      (pll_c2_clk),                                                //               clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                        //             reset.reset
		.stream_in_startofpacket  (pixel_out_buffer_avalon_dc_buffer_source_startofpacket),    //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (pixel_out_buffer_avalon_dc_buffer_source_endofpacket),      //                  .endofpacket
		.stream_in_valid          (pixel_out_buffer_avalon_dc_buffer_source_valid),            //                  .valid
		.stream_in_ready          (pixel_out_buffer_avalon_dc_buffer_source_ready),            //                  .ready
		.stream_in_data           (pixel_out_buffer_avalon_dc_buffer_source_data),             //                  .data
		.slave_read               (mm_interconnect_0_vga_resampler_avalon_rgb_slave_read),     //  avalon_rgb_slave.read
		.slave_readdata           (mm_interconnect_0_vga_resampler_avalon_rgb_slave_readdata), //                  .readdata
		.stream_out_ready         (vga_resampler_avalon_rgb_source_ready),                     // avalon_rgb_source.ready
		.stream_out_startofpacket (vga_resampler_avalon_rgb_source_startofpacket),             //                  .startofpacket
		.stream_out_endofpacket   (vga_resampler_avalon_rgb_source_endofpacket),               //                  .endofpacket
		.stream_out_valid         (vga_resampler_avalon_rgb_source_valid),                     //                  .valid
		.stream_out_data          (vga_resampler_avalon_rgb_source_data)                       //                  .data
	);

	final_soc_vga_scaler vga_scaler (
		.clk                      (pll_c2_clk),                                    //                  clk.clk
		.reset                    (rst_controller_002_reset_out_reset),            //                reset.reset
		.stream_in_startofpacket  (vga_resampler_avalon_rgb_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (vga_resampler_avalon_rgb_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (vga_resampler_avalon_rgb_source_valid),         //                     .valid
		.stream_in_ready          (vga_resampler_avalon_rgb_source_ready),         //                     .ready
		.stream_in_data           (vga_resampler_avalon_rgb_source_data),          //                     .data
		.stream_out_ready         (vga_scaler_avalon_scaler_source_ready),         // avalon_scaler_source.ready
		.stream_out_startofpacket (vga_scaler_avalon_scaler_source_startofpacket), //                     .startofpacket
		.stream_out_endofpacket   (vga_scaler_avalon_scaler_source_endofpacket),   //                     .endofpacket
		.stream_out_valid         (vga_scaler_avalon_scaler_source_valid),         //                     .valid
		.stream_out_data          (vga_scaler_avalon_scaler_source_data),          //                     .data
		.stream_out_channel       (vga_scaler_avalon_scaler_source_channel)        //                     .channel
	);

	final_soc_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                   (clk_clk),                                                     //                                 clk_0_clk.clk
		.PLL_c0_clk                                      (pll_c0_clk),                                                  //                                    PLL_c0.clk
		.PLL_c2_clk                                      (pll_c2_clk),                                                  //                                    PLL_c2.clk
		.GPU_CORE_0_RESET_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                              //    GPU_CORE_0_RESET_reset_bridge_in_reset.reset
		.SDRAM_reset_reset_bridge_in_reset_reset         (rst_controller_001_reset_out_reset),                          //         SDRAM_reset_reset_bridge_in_reset.reset
		.timer_0_reset_reset_bridge_in_reset_reset       (rst_controller_003_reset_out_reset),                          //       timer_0_reset_reset_bridge_in_reset.reset
		.vga_resampler_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                          // vga_resampler_reset_reset_bridge_in_reset.reset
		.GPU_CORE_0_GPU_MASTER_address                   (gpu_core_0_gpu_master_address),                               //                     GPU_CORE_0_GPU_MASTER.address
		.GPU_CORE_0_GPU_MASTER_waitrequest               (gpu_core_0_gpu_master_waitrequest),                           //                                          .waitrequest
		.GPU_CORE_0_GPU_MASTER_chipselect                (gpu_core_0_gpu_master_chipselect),                            //                                          .chipselect
		.GPU_CORE_0_GPU_MASTER_read                      (gpu_core_0_gpu_master_read),                                  //                                          .read
		.GPU_CORE_0_GPU_MASTER_readdata                  (gpu_core_0_gpu_master_readdata),                              //                                          .readdata
		.GPU_CORE_0_GPU_MASTER_readdatavalid             (gpu_core_0_gpu_master_readdatavalid),                         //                                          .readdatavalid
		.GPU_CORE_0_GPU_MASTER_write                     (gpu_core_0_gpu_master_write),                                 //                                          .write
		.GPU_CORE_0_GPU_MASTER_writedata                 (gpu_core_0_gpu_master_writedata),                             //                                          .writedata
		.GPU_CORE_0_GPU_MASTER_response                  (gpu_core_0_gpu_master_response),                              //                                          .response
		.GPU_CORE_0_GPU_MASTER_writeresponsevalid        (gpu_core_0_gpu_master_writeresponsevalid),                    //                                          .writeresponsevalid
		.NIOS2_data_master_address                       (nios2_data_master_address),                                   //                         NIOS2_data_master.address
		.NIOS2_data_master_waitrequest                   (nios2_data_master_waitrequest),                               //                                          .waitrequest
		.NIOS2_data_master_byteenable                    (nios2_data_master_byteenable),                                //                                          .byteenable
		.NIOS2_data_master_read                          (nios2_data_master_read),                                      //                                          .read
		.NIOS2_data_master_readdata                      (nios2_data_master_readdata),                                  //                                          .readdata
		.NIOS2_data_master_write                         (nios2_data_master_write),                                     //                                          .write
		.NIOS2_data_master_writedata                     (nios2_data_master_writedata),                                 //                                          .writedata
		.NIOS2_data_master_debugaccess                   (nios2_data_master_debugaccess),                               //                                          .debugaccess
		.NIOS2_instruction_master_address                (nios2_instruction_master_address),                            //                  NIOS2_instruction_master.address
		.NIOS2_instruction_master_waitrequest            (nios2_instruction_master_waitrequest),                        //                                          .waitrequest
		.NIOS2_instruction_master_read                   (nios2_instruction_master_read),                               //                                          .read
		.NIOS2_instruction_master_readdata               (nios2_instruction_master_readdata),                           //                                          .readdata
		.pixel_dma_avalon_pixel_dma_master_address       (pixel_dma_avalon_pixel_dma_master_address),                   //         pixel_dma_avalon_pixel_dma_master.address
		.pixel_dma_avalon_pixel_dma_master_waitrequest   (pixel_dma_avalon_pixel_dma_master_waitrequest),               //                                          .waitrequest
		.pixel_dma_avalon_pixel_dma_master_read          (pixel_dma_avalon_pixel_dma_master_read),                      //                                          .read
		.pixel_dma_avalon_pixel_dma_master_readdata      (pixel_dma_avalon_pixel_dma_master_readdata),                  //                                          .readdata
		.pixel_dma_avalon_pixel_dma_master_readdatavalid (pixel_dma_avalon_pixel_dma_master_readdatavalid),             //                                          .readdatavalid
		.pixel_dma_avalon_pixel_dma_master_lock          (pixel_dma_avalon_pixel_dma_master_lock),                      //                                          .lock
		.frame_buffer_s1_address                         (mm_interconnect_0_frame_buffer_s1_address),                   //                           frame_buffer_s1.address
		.frame_buffer_s1_write                           (mm_interconnect_0_frame_buffer_s1_write),                     //                                          .write
		.frame_buffer_s1_readdata                        (mm_interconnect_0_frame_buffer_s1_readdata),                  //                                          .readdata
		.frame_buffer_s1_writedata                       (mm_interconnect_0_frame_buffer_s1_writedata),                 //                                          .writedata
		.frame_buffer_s1_byteenable                      (mm_interconnect_0_frame_buffer_s1_byteenable),                //                                          .byteenable
		.frame_buffer_s1_chipselect                      (mm_interconnect_0_frame_buffer_s1_chipselect),                //                                          .chipselect
		.frame_buffer_s1_clken                           (mm_interconnect_0_frame_buffer_s1_clken),                     //                                          .clken
		.frame_buffer_s2_address                         (mm_interconnect_0_frame_buffer_s2_address),                   //                           frame_buffer_s2.address
		.frame_buffer_s2_write                           (mm_interconnect_0_frame_buffer_s2_write),                     //                                          .write
		.frame_buffer_s2_readdata                        (mm_interconnect_0_frame_buffer_s2_readdata),                  //                                          .readdata
		.frame_buffer_s2_writedata                       (mm_interconnect_0_frame_buffer_s2_writedata),                 //                                          .writedata
		.frame_buffer_s2_byteenable                      (mm_interconnect_0_frame_buffer_s2_byteenable),                //                                          .byteenable
		.frame_buffer_s2_chipselect                      (mm_interconnect_0_frame_buffer_s2_chipselect),                //                                          .chipselect
		.frame_buffer_s2_clken                           (mm_interconnect_0_frame_buffer_s2_clken),                     //                                          .clken
		.GPU_CORE_0_GPU_SLAVE_address                    (mm_interconnect_0_gpu_core_0_gpu_slave_address),              //                      GPU_CORE_0_GPU_SLAVE.address
		.GPU_CORE_0_GPU_SLAVE_write                      (mm_interconnect_0_gpu_core_0_gpu_slave_write),                //                                          .write
		.GPU_CORE_0_GPU_SLAVE_read                       (mm_interconnect_0_gpu_core_0_gpu_slave_read),                 //                                          .read
		.GPU_CORE_0_GPU_SLAVE_readdata                   (mm_interconnect_0_gpu_core_0_gpu_slave_readdata),             //                                          .readdata
		.GPU_CORE_0_GPU_SLAVE_writedata                  (mm_interconnect_0_gpu_core_0_gpu_slave_writedata),            //                                          .writedata
		.GPU_CORE_0_GPU_SLAVE_chipselect                 (mm_interconnect_0_gpu_core_0_gpu_slave_chipselect),           //                                          .chipselect
		.jtag_uart_0_avalon_jtag_slave_address           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //             jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                          .write
		.jtag_uart_0_avalon_jtag_slave_read              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                          .read
		.jtag_uart_0_avalon_jtag_slave_readdata          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                          .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                          .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                          .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                          .chipselect
		.keycode_s1_address                              (mm_interconnect_0_keycode_s1_address),                        //                                keycode_s1.address
		.keycode_s1_write                                (mm_interconnect_0_keycode_s1_write),                          //                                          .write
		.keycode_s1_readdata                             (mm_interconnect_0_keycode_s1_readdata),                       //                                          .readdata
		.keycode_s1_writedata                            (mm_interconnect_0_keycode_s1_writedata),                      //                                          .writedata
		.keycode_s1_chipselect                           (mm_interconnect_0_keycode_s1_chipselect),                     //                                          .chipselect
		.NIOS2_debug_mem_slave_address                   (mm_interconnect_0_nios2_debug_mem_slave_address),             //                     NIOS2_debug_mem_slave.address
		.NIOS2_debug_mem_slave_write                     (mm_interconnect_0_nios2_debug_mem_slave_write),               //                                          .write
		.NIOS2_debug_mem_slave_read                      (mm_interconnect_0_nios2_debug_mem_slave_read),                //                                          .read
		.NIOS2_debug_mem_slave_readdata                  (mm_interconnect_0_nios2_debug_mem_slave_readdata),            //                                          .readdata
		.NIOS2_debug_mem_slave_writedata                 (mm_interconnect_0_nios2_debug_mem_slave_writedata),           //                                          .writedata
		.NIOS2_debug_mem_slave_byteenable                (mm_interconnect_0_nios2_debug_mem_slave_byteenable),          //                                          .byteenable
		.NIOS2_debug_mem_slave_waitrequest               (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),         //                                          .waitrequest
		.NIOS2_debug_mem_slave_debugaccess               (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),         //                                          .debugaccess
		.otg_hpi_address_s1_address                      (mm_interconnect_0_otg_hpi_address_s1_address),                //                        otg_hpi_address_s1.address
		.otg_hpi_address_s1_write                        (mm_interconnect_0_otg_hpi_address_s1_write),                  //                                          .write
		.otg_hpi_address_s1_readdata                     (mm_interconnect_0_otg_hpi_address_s1_readdata),               //                                          .readdata
		.otg_hpi_address_s1_writedata                    (mm_interconnect_0_otg_hpi_address_s1_writedata),              //                                          .writedata
		.otg_hpi_address_s1_chipselect                   (mm_interconnect_0_otg_hpi_address_s1_chipselect),             //                                          .chipselect
		.otg_hpi_cs_s1_address                           (mm_interconnect_0_otg_hpi_cs_s1_address),                     //                             otg_hpi_cs_s1.address
		.otg_hpi_cs_s1_write                             (mm_interconnect_0_otg_hpi_cs_s1_write),                       //                                          .write
		.otg_hpi_cs_s1_readdata                          (mm_interconnect_0_otg_hpi_cs_s1_readdata),                    //                                          .readdata
		.otg_hpi_cs_s1_writedata                         (mm_interconnect_0_otg_hpi_cs_s1_writedata),                   //                                          .writedata
		.otg_hpi_cs_s1_chipselect                        (mm_interconnect_0_otg_hpi_cs_s1_chipselect),                  //                                          .chipselect
		.otg_hpi_data_s1_address                         (mm_interconnect_0_otg_hpi_data_s1_address),                   //                           otg_hpi_data_s1.address
		.otg_hpi_data_s1_write                           (mm_interconnect_0_otg_hpi_data_s1_write),                     //                                          .write
		.otg_hpi_data_s1_readdata                        (mm_interconnect_0_otg_hpi_data_s1_readdata),                  //                                          .readdata
		.otg_hpi_data_s1_writedata                       (mm_interconnect_0_otg_hpi_data_s1_writedata),                 //                                          .writedata
		.otg_hpi_data_s1_chipselect                      (mm_interconnect_0_otg_hpi_data_s1_chipselect),                //                                          .chipselect
		.otg_hpi_r_s1_address                            (mm_interconnect_0_otg_hpi_r_s1_address),                      //                              otg_hpi_r_s1.address
		.otg_hpi_r_s1_write                              (mm_interconnect_0_otg_hpi_r_s1_write),                        //                                          .write
		.otg_hpi_r_s1_readdata                           (mm_interconnect_0_otg_hpi_r_s1_readdata),                     //                                          .readdata
		.otg_hpi_r_s1_writedata                          (mm_interconnect_0_otg_hpi_r_s1_writedata),                    //                                          .writedata
		.otg_hpi_r_s1_chipselect                         (mm_interconnect_0_otg_hpi_r_s1_chipselect),                   //                                          .chipselect
		.otg_hpi_reset_s1_address                        (mm_interconnect_0_otg_hpi_reset_s1_address),                  //                          otg_hpi_reset_s1.address
		.otg_hpi_reset_s1_write                          (mm_interconnect_0_otg_hpi_reset_s1_write),                    //                                          .write
		.otg_hpi_reset_s1_readdata                       (mm_interconnect_0_otg_hpi_reset_s1_readdata),                 //                                          .readdata
		.otg_hpi_reset_s1_writedata                      (mm_interconnect_0_otg_hpi_reset_s1_writedata),                //                                          .writedata
		.otg_hpi_reset_s1_chipselect                     (mm_interconnect_0_otg_hpi_reset_s1_chipselect),               //                                          .chipselect
		.otg_hpi_w_s1_address                            (mm_interconnect_0_otg_hpi_w_s1_address),                      //                              otg_hpi_w_s1.address
		.otg_hpi_w_s1_write                              (mm_interconnect_0_otg_hpi_w_s1_write),                        //                                          .write
		.otg_hpi_w_s1_readdata                           (mm_interconnect_0_otg_hpi_w_s1_readdata),                     //                                          .readdata
		.otg_hpi_w_s1_writedata                          (mm_interconnect_0_otg_hpi_w_s1_writedata),                    //                                          .writedata
		.otg_hpi_w_s1_chipselect                         (mm_interconnect_0_otg_hpi_w_s1_chipselect),                   //                                          .chipselect
		.pixel_dma_avalon_control_slave_address          (mm_interconnect_0_pixel_dma_avalon_control_slave_address),    //            pixel_dma_avalon_control_slave.address
		.pixel_dma_avalon_control_slave_write            (mm_interconnect_0_pixel_dma_avalon_control_slave_write),      //                                          .write
		.pixel_dma_avalon_control_slave_read             (mm_interconnect_0_pixel_dma_avalon_control_slave_read),       //                                          .read
		.pixel_dma_avalon_control_slave_readdata         (mm_interconnect_0_pixel_dma_avalon_control_slave_readdata),   //                                          .readdata
		.pixel_dma_avalon_control_slave_writedata        (mm_interconnect_0_pixel_dma_avalon_control_slave_writedata),  //                                          .writedata
		.pixel_dma_avalon_control_slave_byteenable       (mm_interconnect_0_pixel_dma_avalon_control_slave_byteenable), //                                          .byteenable
		.PLL_pll_slave_address                           (mm_interconnect_0_pll_pll_slave_address),                     //                             PLL_pll_slave.address
		.PLL_pll_slave_write                             (mm_interconnect_0_pll_pll_slave_write),                       //                                          .write
		.PLL_pll_slave_read                              (mm_interconnect_0_pll_pll_slave_read),                        //                                          .read
		.PLL_pll_slave_readdata                          (mm_interconnect_0_pll_pll_slave_readdata),                    //                                          .readdata
		.PLL_pll_slave_writedata                         (mm_interconnect_0_pll_pll_slave_writedata),                   //                                          .writedata
		.SDRAM_s1_address                                (mm_interconnect_0_sdram_s1_address),                          //                                  SDRAM_s1.address
		.SDRAM_s1_write                                  (mm_interconnect_0_sdram_s1_write),                            //                                          .write
		.SDRAM_s1_read                                   (mm_interconnect_0_sdram_s1_read),                             //                                          .read
		.SDRAM_s1_readdata                               (mm_interconnect_0_sdram_s1_readdata),                         //                                          .readdata
		.SDRAM_s1_writedata                              (mm_interconnect_0_sdram_s1_writedata),                        //                                          .writedata
		.SDRAM_s1_byteenable                             (mm_interconnect_0_sdram_s1_byteenable),                       //                                          .byteenable
		.SDRAM_s1_readdatavalid                          (mm_interconnect_0_sdram_s1_readdatavalid),                    //                                          .readdatavalid
		.SDRAM_s1_waitrequest                            (mm_interconnect_0_sdram_s1_waitrequest),                      //                                          .waitrequest
		.SDRAM_s1_chipselect                             (mm_interconnect_0_sdram_s1_chipselect),                       //                                          .chipselect
		.timer_0_s1_address                              (mm_interconnect_0_timer_0_s1_address),                        //                                timer_0_s1.address
		.timer_0_s1_write                                (mm_interconnect_0_timer_0_s1_write),                          //                                          .write
		.timer_0_s1_readdata                             (mm_interconnect_0_timer_0_s1_readdata),                       //                                          .readdata
		.timer_0_s1_writedata                            (mm_interconnect_0_timer_0_s1_writedata),                      //                                          .writedata
		.timer_0_s1_chipselect                           (mm_interconnect_0_timer_0_s1_chipselect),                     //                                          .chipselect
		.vga_resampler_avalon_rgb_slave_read             (mm_interconnect_0_vga_resampler_avalon_rgb_slave_read),       //            vga_resampler_avalon_rgb_slave.read
		.vga_resampler_avalon_rgb_slave_readdata         (mm_interconnect_0_vga_resampler_avalon_rgb_slave_readdata)    //                                          .readdata
	);

	final_soc_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_irq_irq)                   //    sender.irq
	);

	final_soc_avalon_st_adapter #(
		.inBitsPerSymbol (10),
		.inUsePackets    (1),
		.inDataWidth     (30),
		.inChannelWidth  (2),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (30),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (pll_c2_clk),                                    // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_002_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (vga_scaler_avalon_scaler_source_data),          //     in_0.data
		.in_0_valid          (vga_scaler_avalon_scaler_source_valid),         //         .valid
		.in_0_ready          (vga_scaler_avalon_scaler_source_ready),         //         .ready
		.in_0_startofpacket  (vga_scaler_avalon_scaler_source_startofpacket), //         .startofpacket
		.in_0_endofpacket    (vga_scaler_avalon_scaler_source_endofpacket),   //         .endofpacket
		.in_0_channel        (vga_scaler_avalon_scaler_source_channel),       //         .channel
		.out_0_data          (avalon_st_adapter_out_0_data),                  //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),                 //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),                 //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),         //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket)            //         .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios2_debug_reset_request_reset),    // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios2_debug_reset_request_reset),    // reset_in1.reset
		.clk            (pll_c0_clk),                         //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios2_debug_reset_request_reset),    // reset_in1.reset
		.clk            (pll_c2_clk),                         //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
